`ifndef CONV_CONFIGURATION_PKG_SV
    `define CONV_CONFIGURATION_PKG_SV


package conv_configuration_pkg;


    // Include uvm package and uvm macros and config file        
     import uvm_pkg::*;     
    `include "uvm_macros.svh" 
    `include "conv_config.sv" 


endpackage : conv_configuration_pkg


`endif   